** Profile: "SCHEMATIC1-sim"  [ E:\DOCTORADO\MiniCycling\Modelado_planta\5-TrabajoPandemia\7-TestDelModeloPID\OBT\4-Analisis de fallas por desviacion\Analisis de fallas no detectadas\9a-ModeloOrcad_conPID_STD18\fuentermnconpid-pspicefiles\schematic1\sim.sim ] 

** Creating circuit file "sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\delfi\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "C:\Cadence\SPB_16.6\tools\pspice\library\AD8170.lib" 
.lib "C:\Cadence\SPB_16.6\tools\pspice\library\LMH7324.lib" 
.lib "C:\Cadence\SPB_16.6\tools\pspice\library\IXTN660N04T4.lib" 
.lib "C:\Cadence\SPB_16.6\tools\pspice\library\t5kp10a.lib" 
.lib "C:\Cadence\SPB_16.6\tools\pspice\library\MAX4376H.lib" 
.lib "C:\Cadence\SPB_16.6\tools\pspice\library\STD18NF03Lmodif.lib" 
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 100us 0 10n 
.STEP PARAM cap LIST 235p, 470p, 705p 
.OPTIONS ADVCONV
.OPTIONS ABSTOL= 10.0p
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
